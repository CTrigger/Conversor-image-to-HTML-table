0 => (0 => (0,0,15), 1 => (0,0,15), 2 => (0,0,15), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (0,0,15), 8 => (0,0,15), 9 => (0,0,15)), 
1 => (0 => (0,0,15), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (0,0,15)), 
2 => (0 => (0,0,15), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (0,0,15)), 
3 => (0 => (15,15,0), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (15,15,0)), 
4 => (0 => (15,15,0), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (15,15,0)), 
5 => (0 => (15,15,0), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (15,15,0)), 
6 => (0 => (15,15,0), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (0,0,15), 5 => (0,0,15), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (15,15,0)), 
7 => (0 => (0,0,15), 1 => (15,15,0), 2 => (15,15,0), 3 => (0,0,15), 4 => (0,0,15), 5 => (0,0,15), 6 => (0,0,15), 7 => (15,15,0), 8 => (15,15,0), 9 => (0,0,15)), 
8 => (0 => (0,0,15), 1 => (15,15,0), 2 => (0,0,15), 3 => (0,0,15), 4 => (0,0,15), 5 => (0,0,15), 6 => (0,0,15), 7 => (0,0,15), 8 => (15,15,0), 9 => (0,0,15)), 
9 => (0 => (0,0,15), 1 => (0,0,15), 2 => (0,0,15), 3 => (0,0,15), 4 => (0,0,15), 5 => (0,0,15), 6 => (0,0,15), 7 => (0,0,15), 8 => (0,0,15), 9 => (0,0,15)) 
